`timescale 1ns / 1ps

module test(

    );
	reg ACLK, ARESETN;
    reg [31:0]S_AXIS_TDATA;
    reg S_AXIS_TVALID, M_AXIS_TREADY, S_AXIS_TLAST;
    wire [31:0]M_AXIS_TDATA;
    wire M_AXIS_TVALID, S_AXIS_TREADY;

    myip_v1_0 dut(ACLK,
        ARESETN,
        S_AXIS_TREADY,
        S_AXIS_TDATA,
        S_AXIS_TLAST,
        S_AXIS_TVALID,
        M_AXIS_TVALID,
        M_AXIS_TDATA,
        M_AXIS_TLAST,
        M_AXIS_TREADY);

    reg i;
    initial begin
        ACLK = 0;
        i = 0;
        #3;
        ARESETN = 0;
        #20; 
        ARESETN = 1; 
        M_AXIS_TREADY = 1;
        #10;
        S_AXIS_TVALID = 1;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd216;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd224;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd52;
        #10;
        S_AXIS_TDATA = 32'd40;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd212;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd208;
        #10;
        S_AXIS_TDATA = 32'd200;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd196;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd204;
        #10;
        S_AXIS_TDATA = 32'd220;
        #10;
        S_AXIS_TDATA = 32'd128;
        #10;
        S_AXIS_TDATA = 32'd228;
        #10;
        S_AXIS_TDATA = 32'd192;
        #10;
        S_AXIS_TDATA = 32'd4294966608;
        #10;
        S_AXIS_TDATA = 32'd4294967233;
        #10;
        S_AXIS_TDATA = 32'd4294966280;
        #10;
        S_AXIS_TDATA = 32'd4294965672;
        #10;
        S_AXIS_TDATA = 32'd4294961584;
        #10;
        S_AXIS_TDATA = 32'd4294966108;
        #10;
        S_AXIS_TDATA = 32'd4294966771;
        #10;
        S_AXIS_TDATA = 32'd4294966579;
        #10;
        S_AXIS_TDATA = 32'd4294965888;
        #10;
        S_AXIS_TDATA = 32'd4294965571;
        #10;
        S_AXIS_TDATA = 32'd4294966995;
        #10;
        S_AXIS_TDATA = 32'd4294967060;
        #10;
        S_AXIS_TDATA = 32'd4294966803;
        #10;
        S_AXIS_TDATA = 32'd4294966260;
        #10;
        S_AXIS_TDATA = 32'd4294966881;
        #10;
        S_AXIS_TDATA = 32'd4294966495;
        #10;
        S_AXIS_TDATA = 32'd4294967190;
        #10;
        S_AXIS_TDATA = 32'd4294966534;
        #10;
        S_AXIS_TDATA = 32'd4294967033;
        #10;
        S_AXIS_TDATA = 32'd4294966361;
        #10;
        S_AXIS_TDATA = 32'd4294967007;
        #10;
        S_AXIS_TDATA = 32'd4294967272;
        #10;
        S_AXIS_TDATA = 32'd54;
        #10;
        S_AXIS_TDATA = 32'd4294966520;
        #10;
        S_AXIS_TDATA = 32'd4294966947;
        #10;
        S_AXIS_TDATA = 32'd4294966592;
        #10;
        S_AXIS_TDATA = 32'd490;
        #10;
        S_AXIS_TDATA = 32'd37;
        #10;
        S_AXIS_TDATA = 32'd133;
        #10;
        S_AXIS_TDATA = 32'd4294965650;
        #10;
        S_AXIS_TDATA = 32'd4294966111;
        #10;
        S_AXIS_TDATA = 32'd521;
        #10;
        S_AXIS_TDATA = 32'd472;
        #10;
        S_AXIS_TDATA = 32'd111;
        #10;
        S_AXIS_TDATA = 32'd4294966464;
        #10;
        S_AXIS_TDATA = 32'd4294965705;
        #10;
        S_AXIS_TDATA = 32'd4971;
        #10;
        S_AXIS_TDATA = 32'd715;
        #10;
        S_AXIS_TDATA = 32'd4325;
        #10;
        S_AXIS_TDATA = 32'd602;
        #10;
        S_AXIS_TDATA = 32'd119;
        #10;
        S_AXIS_TDATA = 32'd4294966090;
        #10;
        S_AXIS_TDATA = 32'd4294959058;
        #10;
        S_AXIS_TDATA = 32'd421;
        #10;
        S_AXIS_TDATA = 32'd4294963351;
        #10;
        S_AXIS_TDATA = 32'd2148;
        #10;
        S_AXIS_TDATA = 32'd4294961017;
        #10;
        S_AXIS_TDATA = 32'd4294961720;
        #10;
        S_AXIS_TDATA = 32'd2270;
        #10;
        S_AXIS_TDATA = 32'd820;
        #10;
        S_AXIS_TDATA = 32'd694;
        #10;
        S_AXIS_TDATA = 32'd4294967051;
        #10;
        S_AXIS_TDATA = 32'd780;
        #10;
        S_AXIS_TDATA = 32'd4294967144;
        #10;
        S_AXIS_TDATA = 32'd4294967163;
        #10;
        S_AXIS_TDATA = 32'd4294965205;
        #10;
        S_AXIS_TDATA = 32'd4294966569;
        #10;
        S_AXIS_TDATA = 32'd4294965811;
        #10;
        S_AXIS_TDATA = 32'd565;
        #10;
        S_AXIS_TDATA = 32'd4294966214;
        #10;
        S_AXIS_TDATA = 32'd4294966734;
        #10;
        S_AXIS_TDATA = 32'd4294966126;
        #10;
        S_AXIS_TDATA = 32'd7434;
        #10;
        S_AXIS_TDATA = 32'd1040;
        #10;
        S_AXIS_TDATA = 32'd4504;
        #10;
        S_AXIS_TDATA = 32'd4294962458;
        #10;
        S_AXIS_TDATA = 32'd1737;
        #10;
        S_AXIS_TDATA = 32'd4294965967;
        #10;
        S_AXIS_TDATA = 32'd2465;
        #10;
        S_AXIS_TDATA = 32'd791;
        #10;
        S_AXIS_TDATA = 32'd4294965583;
        #10;
        S_AXIS_TDATA = 32'd2100;
        #10;
        S_AXIS_TDATA = 32'd4294960669;
        #10;
        S_AXIS_TDATA = 32'd218;
        #10;
        S_AXIS_TDATA = 32'd7914;
        #10;
        S_AXIS_TDATA = 32'd1698;
        #10;
        S_AXIS_TDATA = 32'd935;
        #10;
        S_AXIS_TDATA = 32'd849;
        #10;
        S_AXIS_TDATA = 32'd4294965804;
        #10;
        S_AXIS_TDATA = 32'd382;
        #10;
        S_AXIS_TDATA = 32'd4294966221;
        #10;
        S_AXIS_TDATA = 32'd1278;
        #10;
        S_AXIS_TDATA = 32'd4294967007;
        #10;
        S_AXIS_TDATA = 32'd4294966023;
        #10;
        S_AXIS_TDATA = 32'd599;
        #10;
        S_AXIS_TDATA = 32'd4294966370;
        #10;
        S_AXIS_TDATA = 32'd75;
        #10;
        S_AXIS_TDATA = 32'd1967;
        #10;
        S_AXIS_TDATA = 32'd368;
        #10;
        S_AXIS_TDATA = 32'd4294966876;
        #10;
        S_AXIS_TDATA = 32'd4294967212;
        #10;
        S_AXIS_TDATA = 32'd722;
        #10;
        S_AXIS_TDATA = 32'd4294966247;
        #10;
        S_AXIS_TDATA = 32'd84;
        #10;
        S_AXIS_TDATA = 32'd4294966028;
        #10;
        S_AXIS_TDATA = 32'd4294965977;
        #10;
        S_AXIS_TDATA = 32'd4294966969;
        #10;
        S_AXIS_TDATA = 32'd381;
        #10;
        S_AXIS_TDATA = 32'd4294966315;
        #10;
        S_AXIS_TDATA = 32'd4294966979;
        #10;
        S_AXIS_TDATA = 32'd4294965798;
        #10;
        S_AXIS_TDATA = 32'd4294967171;
        #10;
        S_AXIS_TDATA = 32'd54;
        #10;
        S_AXIS_TDATA = 32'd4294967093;
        #10;
        S_AXIS_TDATA = 32'd334;
        #10;
        S_AXIS_TDATA = 32'd4294967027;
        #10;
        S_AXIS_TDATA = 32'd4294966533;
        #10;
        S_AXIS_TDATA = 32'd4294966022;
        #10;
        S_AXIS_TDATA = 32'd334;
        #10;
        S_AXIS_TDATA = 32'd4294966379;
        #10;
        S_AXIS_TDATA = 32'd394;
        #10;
        S_AXIS_TDATA = 32'd4294966350;
        #10;
        S_AXIS_TDATA = 32'd4294966145;
        #10;
        S_AXIS_TDATA = 32'd4294966991;
        #10;
        S_AXIS_TDATA = 32'd847;
        #10;
        S_AXIS_TDATA = 32'd126;
        #10;
        S_AXIS_TDATA = 32'd185;
        #10;
        S_AXIS_TDATA = 32'd4294965666;
        #10;
        S_AXIS_TDATA = 32'd67;
        #10;
        S_AXIS_TDATA = 32'd4294966206;
        #10;
        S_AXIS_TDATA = 32'd811;
        #10;
        S_AXIS_TDATA = 32'd289;
        #10;
        S_AXIS_TDATA = 32'd4294966318;
        #10;
        S_AXIS_TDATA = 32'd4294966647;
        #10;
        S_AXIS_TDATA = 32'd4294966341;
        #10;
        S_AXIS_TDATA = 32'd4294967179;
        #10;
        S_AXIS_TDATA = 32'd923;
        #10;
        S_AXIS_TDATA = 32'd4294966750;
        #10;
        S_AXIS_TDATA = 32'd4294965074;
        #10;
        S_AXIS_TDATA = 32'd214;
        #10;
        S_AXIS_TDATA = 32'd4294967051;
        #10;
        S_AXIS_TDATA = 32'd736;
        #10;
        S_AXIS_TDATA = 32'd4294967166;
        #10;
        S_AXIS_TDATA = 32'd313;
        #10;
        S_AXIS_TDATA = 32'd4294966132;
        #10;
        S_AXIS_TDATA = 32'd2451;
        #10;
        S_AXIS_TDATA = 32'd4294967156;
        #10;
        S_AXIS_TDATA = 32'd4294966683;
        #10;
        S_AXIS_TDATA = 32'd4294966070;
        #10;
        S_AXIS_TDATA = 32'd36;
        #10;
        S_AXIS_TDATA = 32'd698;
        #10;
        S_AXIS_TDATA = 32'd4294966779;
        #10;
        S_AXIS_TDATA = 32'd4294966270;
        #10;
        S_AXIS_TDATA = 32'd9249;
        #10;
        S_AXIS_TDATA = 32'd1055;
        #10;
        S_AXIS_TDATA = 32'd4294965436;
        #10;
        S_AXIS_TDATA = 32'd440;
        #10;
        S_AXIS_TDATA = 32'd373;
        #10;
        S_AXIS_TDATA = 32'd4294966773;
        #10;
        S_AXIS_TDATA = 32'd88;
        #10;
        S_AXIS_TDATA = 32'd722;
        #10
        S_AXIS_TVALID = 0;
        S_AXIS_TDATA = 0;
    end

    always begin
    	#5; ACLK = ~ACLK;
    end
        
        
endmodule
